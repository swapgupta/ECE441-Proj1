library verilog;
use verilog.vl_types.all;
entity proj1_tb is
end proj1_tb;
