library verilog;
use verilog.vl_types.all;
entity parity_tb is
end parity_tb;
